Wire declaration;

`default_nettype none
module top_module(
    input a,
    input b,
    input c,
    input d,
    output out,
    output out_n   ); 
    wire ab , cd;
    assign ab = a & b;
    assign cd = c & d;
    assign out = ab | cd;
    assign out_n = ~(ab | cd);

endmodule

7458;

module top_module ( 
    input p1a, p1b, p1c, p1d, p1e, p1f,
    output p1y,
    input p2a, p2b, p2c, p2d,
    output p2y );
    assign p1y = (p1a & p1b & p1c) | (p1d & p1e & p1f);
    assign p2y = (p2a & p2b) | (p2c & p2d);


endmodule